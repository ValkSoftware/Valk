module util

import time

__global uptime = time.new_stopwatch()