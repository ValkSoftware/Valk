module chat

enum TextStyle {
	bold
	under
	strike
	obfusc
	italic
	normal
}

